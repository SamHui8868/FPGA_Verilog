library verilog;
use verilog.vl_types.all;
entity fDIV25K_vlg_vec_tst is
end fDIV25K_vlg_vec_tst;
