library verilog;
use verilog.vl_types.all;
entity hw5_vlg_vec_tst is
end hw5_vlg_vec_tst;
