library verilog;
use verilog.vl_types.all;
entity fDIV27M_vlg_vec_tst is
end fDIV27M_vlg_vec_tst;
