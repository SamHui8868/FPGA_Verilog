library verilog;
use verilog.vl_types.all;
entity serial_out_vlg_vec_tst is
end serial_out_vlg_vec_tst;
