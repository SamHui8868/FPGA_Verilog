library verilog;
use verilog.vl_types.all;
entity TPC_vlg_vec_tst is
end TPC_vlg_vec_tst;
