library verilog;
use verilog.vl_types.all;
entity hw2_vlg_check_tst is
    port(
        \_A\            : in     vl_logic;
        \_B\            : in     vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end hw2_vlg_check_tst;
