library verilog;
use verilog.vl_types.all;
entity stepMotorctr_vlg_vec_tst is
end stepMotorctr_vlg_vec_tst;
