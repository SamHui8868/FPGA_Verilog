library verilog;
use verilog.vl_types.all;
entity FDIV50K_vlg_vec_tst is
end FDIV50K_vlg_vec_tst;
