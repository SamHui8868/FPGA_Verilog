library verilog;
use verilog.vl_types.all;
entity SO_vlg_check_tst is
    port(
        dout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end SO_vlg_check_tst;
