library verilog;
use verilog.vl_types.all;
entity Fdiv_Beat_vlg_check_tst is
    port(
        Fout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Fdiv_Beat_vlg_check_tst;
