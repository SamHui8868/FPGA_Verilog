library verilog;
use verilog.vl_types.all;
entity Comparator_vlg_vec_tst is
end Comparator_vlg_vec_tst;
