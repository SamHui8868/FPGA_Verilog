library verilog;
use verilog.vl_types.all;
entity FDIV50K is
    port(
        fin             : in     vl_logic;
        fout            : out    vl_logic
    );
end FDIV50K;
