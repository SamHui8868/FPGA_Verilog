library verilog;
use verilog.vl_types.all;
entity FDIV25K_vlg_vec_tst is
end FDIV25K_vlg_vec_tst;
