library verilog;
use verilog.vl_types.all;
entity serial_out_vlg_check_tst is
    port(
        D               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end serial_out_vlg_check_tst;
