library verilog;
use verilog.vl_types.all;
entity fDIV27M_vlg_check_tst is
    port(
        fout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fDIV27M_vlg_check_tst;
