library verilog;
use verilog.vl_types.all;
entity \_output_vlg_check_tst\ is
    port(
        reset           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end \_output_vlg_check_tst\;
