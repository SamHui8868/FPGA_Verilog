library verilog;
use verilog.vl_types.all;
entity Mux2to1_5_vlg_vec_tst is
end Mux2to1_5_vlg_vec_tst;
