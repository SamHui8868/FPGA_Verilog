library verilog;
use verilog.vl_types.all;
entity hw4_vlg_vec_tst is
end hw4_vlg_vec_tst;
