library verilog;
use verilog.vl_types.all;
entity AGU_vlg_vec_tst is
end AGU_vlg_vec_tst;
