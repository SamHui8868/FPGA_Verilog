library verilog;
use verilog.vl_types.all;
entity Asyn_counter_vlg_vec_tst is
end Asyn_counter_vlg_vec_tst;
