library verilog;
use verilog.vl_types.all;
entity hw4_vlg_check_tst is
    port(
        CP              : in     vl_logic;
        D               : in     vl_logic;
        str             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end hw4_vlg_check_tst;
