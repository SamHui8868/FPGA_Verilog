library verilog;
use verilog.vl_types.all;
entity hw4n_vlg_vec_tst is
end hw4n_vlg_vec_tst;
