module ctrl(din,clk,start,str);
input din,clk;
output reg start,str;
reg[1:0]cs,ns;
reg[3:0]count;
always@(posedge din or posedge clk)
start=din;

always@(posedge clk)
cs<=ns;
always@(posedge clk)
case(cs)
2'd0:str<=1'd0;
2'd1:str<=1'd0;
2'd2:str<=1'd0;
2'd3:str<=1'd1;
endcase

always@(posedge clk)
if(cs==2'd2)
count=count+1;
else
count=4'd0;

always@(cs)
case(cs)
2'd0:ns<=(start)?2'd1:2'd0;
2'd1:ns<=2'd2;
2'd2:ns<=(count==4'd14)?2'd3:2'd2;
2'd3:ns<=2'd0;
endcase
endmodule
