library verilog;
use verilog.vl_types.all;
entity Fdiv_Sound_vlg_vec_tst is
end Fdiv_Sound_vlg_vec_tst;
