library verilog;
use verilog.vl_types.all;
entity LEDENC_vlg_vec_tst is
end LEDENC_vlg_vec_tst;
