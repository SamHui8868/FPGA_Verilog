library verilog;
use verilog.vl_types.all;
entity ADctrl_vlg_vec_tst is
end ADctrl_vlg_vec_tst;
