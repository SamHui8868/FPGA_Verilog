library verilog;
use verilog.vl_types.all;
entity FDIV_vlg_vec_tst is
end FDIV_vlg_vec_tst;
