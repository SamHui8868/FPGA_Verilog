library verilog;
use verilog.vl_types.all;
entity hw7_vlg_vec_tst is
end hw7_vlg_vec_tst;
