library verilog;
use verilog.vl_types.all;
entity fDIV27M is
    port(
        fin             : in     vl_logic;
        fout            : out    vl_logic
    );
end fDIV27M;
