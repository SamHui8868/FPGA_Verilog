library verilog;
use verilog.vl_types.all;
entity ADdff8_vlg_vec_tst is
end ADdff8_vlg_vec_tst;
