library verilog;
use verilog.vl_types.all;
entity Dff8_vlg_vec_tst is
end Dff8_vlg_vec_tst;
