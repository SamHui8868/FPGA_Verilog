library verilog;
use verilog.vl_types.all;
entity hw2_vlg_vec_tst is
end hw2_vlg_vec_tst;
