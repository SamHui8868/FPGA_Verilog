library verilog;
use verilog.vl_types.all;
entity \_7segENC_vlg_check_tst\ is
    port(
        \_7seg\         : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end \_7segENC_vlg_check_tst\;
