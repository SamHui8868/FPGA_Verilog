library verilog;
use verilog.vl_types.all;
entity \_output_vlg_vec_tst\ is
end \_output_vlg_vec_tst\;
