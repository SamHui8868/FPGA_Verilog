library verilog;
use verilog.vl_types.all;
entity ADctr_vlg_vec_tst is
end ADctr_vlg_vec_tst;
