module ADdff8(clk,en,din,dout);
input clk,en;
input [7:0]din;
output reg[7:0]dout;
always @(posedge clk)
dout=(en==1'd1)?din:dout;
endmodule	