library verilog;
use verilog.vl_types.all;
entity hw1_vlg_vec_tst is
end hw1_vlg_vec_tst;
