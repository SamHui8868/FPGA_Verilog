library verilog;
use verilog.vl_types.all;
entity ctrl_vlg_vec_tst is
end ctrl_vlg_vec_tst;
