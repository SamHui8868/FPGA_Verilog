library verilog;
use verilog.vl_types.all;
entity Fdiv_Beat_vlg_sample_tst is
    port(
        Fin             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Fdiv_Beat_vlg_sample_tst;
