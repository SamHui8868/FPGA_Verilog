library verilog;
use verilog.vl_types.all;
entity SO_vlg_vec_tst is
end SO_vlg_vec_tst;
