library verilog;
use verilog.vl_types.all;
entity oneshot_vlg_vec_tst is
end oneshot_vlg_vec_tst;
