library verilog;
use verilog.vl_types.all;
entity fDIV50M_vlg_vec_tst is
end fDIV50M_vlg_vec_tst;
