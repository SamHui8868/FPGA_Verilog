library verilog;
use verilog.vl_types.all;
entity fDIV25K_vlg_check_tst is
    port(
        fout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fDIV25K_vlg_check_tst;
