library verilog;
use verilog.vl_types.all;
entity stepMotorctr_vlg_check_tst is
    port(
        smctr           : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end stepMotorctr_vlg_check_tst;
