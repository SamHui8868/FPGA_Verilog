library verilog;
use verilog.vl_types.all;
entity \_7segENC_vlg_vec_tst\ is
end \_7segENC_vlg_vec_tst\;
