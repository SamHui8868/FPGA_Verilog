library verilog;
use verilog.vl_types.all;
entity Fdiv_Beat_vlg_vec_tst is
end Fdiv_Beat_vlg_vec_tst;
