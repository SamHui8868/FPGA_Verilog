library verilog;
use verilog.vl_types.all;
entity sel_DIVN_vlg_vec_tst is
end sel_DIVN_vlg_vec_tst;
