library verilog;
use verilog.vl_types.all;
entity Fdiv_Beat is
    port(
        Fin             : in     vl_logic;
        Fout            : out    vl_logic
    );
end Fdiv_Beat;
