library verilog;
use verilog.vl_types.all;
entity FDIV50K_vlg_check_tst is
    port(
        fout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FDIV50K_vlg_check_tst;
